LIBRARY IEEE; 
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY vhdl IS 
PORT (
		HEX00 : OUT STD_LOGIC;
		HEX01 : OUT STD_LOGIC;
		HEX02 : OUT STD_LOGIC;
		HEX03 : OUT STD_LOGIC;
		HEX04 : OUT STD_LOGIC;
		HEX05 : OUT STD_LOGIC;
		HEX06 : OUT STD_LOGIC;
		HEX10 : OUT STD_LOGIC;
		HEX11 : OUT STD_LOGIC;
		HEX12 : OUT STD_LOGIC;
		HEX13 : OUT STD_LOGIC;
		HEX14 : OUT STD_LOGIC;
		HEX15 : OUT STD_LOGIC;
		HEX16 : OUT STD_LOGIC;
		HEX20 : OUT STD_LOGIC;
		HEX21 : OUT STD_LOGIC;
		HEX22 : OUT STD_LOGIC;
		HEX23 : OUT STD_LOGIC;
		HEX24 : OUT STD_LOGIC;
		HEX25 : OUT STD_LOGIC;
		HEX26 : OUT STD_LOGIC;
		HEX30 : OUT STD_LOGIC;
		HEX31 : OUT STD_LOGIC;
		HEX32 : OUT STD_LOGIC;
		HEX33 : OUT STD_LOGIC;
		HEX34 : OUT STD_LOGIC;
		HEX35 : OUT STD_LOGIC;
		HEX36 : OUT STD_LOGIC;
		HEX40 : OUT STD_LOGIC;
		HEX41 : OUT STD_LOGIC;
		HEX42 : OUT STD_LOGIC;
		HEX43 : OUT STD_LOGIC;
		HEX44 : OUT STD_LOGIC;
		HEX45 : OUT STD_LOGIC;
		HEX46 : OUT STD_LOGIC;
		HEX50 : OUT STD_LOGIC;
		HEX51 : OUT STD_LOGIC;
		HEX52 : OUT STD_LOGIC;
		HEX53 : OUT STD_LOGIC;
		HEX54 : OUT STD_LOGIC;
		HEX55 : OUT STD_LOGIC;
		HEX56 : OUT STD_LOGIC;
		clk: IN STD_LOGIC;
		sw1 : IN STD_LOGIC;
		SW0 : IN STD_LOGIC;
clock_1Hz : OUT STD_LOGIC
		);	
END vhdl;



architecture behavioral of vhdl is
signal i : std_logic_vector(4 downto 0):="00000";
SIGNAL count_1hz : STD_LOGIC_VECTOR(25 DOWNTO 0):= "00000000000000000000000000" ;
SIGNAL  clock_1Hz_int : STD_LOGIC;
BEGIN
PROCESS 
BEGIN

WAIT UNTIL clk'EVENT and clk = '1' ;
IF count_1hz < 9000000 THEN
count_1hz <= count_1hz + 1;
ELSE
count_1hz <= "00000000000000000000000000" ;
END IF;
IF count_1hz < 9000000 THEN
clock_1Hz_int <= '0';
ELSE
clock_1Hz_int <= '1' ;
END IF; 

END PROCESS; 



process(clock_1Hz_int)
begin 
if(rising_edge (clock_1Hz_int) ) 
then 

	

 
if(SW0='1') then
		case i is  
		when "00000" => 
								--cas 1	
	  HEX00 <= '0';
	  HEX01 <= '1';
	  HEX02 <= '0';
	  HEX03 <= '0';
	  HEX04 <= '0';
	  HEX05 <= '0';
	  HEX06 <= '1';
HEX10<='1';
HEX11<='1';
HEX12<='1';
HEX13<='1';
HEX14<='1';
HEX15<='1';
HEX16<='1';
			HEX20<='1';
			HEX21<='1';
			HEX22<='1';
			HEX23<='1';
			HEX24<='1';
			HEX25<='1';
			HEX26<='1';
HEX30<='1';
HEX31<='1';
HEX32<='1';
HEX33<='1';
HEX34<='1';
HEX35<='1';
HEX36<='1';	
		HEX40<='1';
		HEX41<='1';
		HEX42<='1';
		HEX43<='1';
		HEX44<='1';
		HEX45<='1';
		HEX46<='1';
HEX50<='1';
HEX51<='1';
HEX52<='1';
HEX53<='1';
HEX54<='1';
HEX55<='1';
HEX56<='1';
	
	  
	  i <= "00001";
	  
								--cas 2
	  when "00001" => 
	  HEX00<='1';
	  HEX01<='0';
	  HEX02<='0';
	  HEX03<='0';
	  HEX04<='0';
	  HEX05<='0';
	  HEX06<='1' ;
HEX10<='0' ;
HEX11<='1' ;
HEX12<='0' ;
HEX13<='0' ;
HEX14<='0' ;
HEX15<='0' ;
HEX16<='1' ;
		HEX20<='1';
		HEX21<='1';
		HEX22<='1';
		HEX23<='1';
		HEX24<='1';
		HEX25<='1';
		HEX26<='1';
HEX30<='1';
HEX31<='1';
HEX32<='1';
HEX33<='1';
HEX34<='1';
HEX35<='1';
HEX36<='1';
		HEX40<='1';
		HEX41<='1';
		HEX42<='1';
		HEX43<='1';
		HEX44<='1';
		HEX45<='1';
		HEX46<='1';
HEX50<='1';
HEX51<='1';
HEX52<='1';
HEX53<='1';
HEX54<='1';
HEX55<='1';
HEX56<='1';
		

	  i<="00010";
								--cas 3
	  when "00010" => 
	  HEX00<='1';
	  HEX01<='1';
	  HEX02<='1';
	  HEX03<='1';
	  HEX04<='0';
	  HEX05<='0';
	  HEX06<='1' ;
HEX10<='1' ; 
HEX11<='0' ; 
HEX12<='0' ; 
HEX13<='0' ; 
HEX14<='0' ; 
HEX15<='0' ; 
HEX16<='1' ;
		HEX20<='0' ;
		HEX21<='1' ;
		HEX22<='0' ;
		HEX23<='0' ;
		HEX24<='0' ;
		HEX25<='0' ;
		HEX26<='1' ;
HEX30<='1';
HEX31<='1';
HEX32<='1';
HEX33<='1';
HEX34<='1';
HEX35<='1';
HEX36<='1';
		HEX40<='1';
		HEX41<='1';
		HEX42<='1';
		HEX43<='1';
		HEX44<='1';
		HEX45<='1';
		HEX46<='1';
HEX50<='1';
HEX51<='1';
HEX52<='1';
HEX53<='1';
HEX54<='1';
HEX55<='1';
HEX56<='1';
		
	  i<="00011";
							--cas 4
	  when "00011" => 
	  HEX00<='1';
	  HEX01<='1';
	  HEX02<='1';
	  HEX03<='0';
	  HEX04<='0';
	  HEX05<='0';
	  HEX06<='1' ;
HEX10<='1' ; 
HEX11<='1' ; 
HEX12<='1' ; 
HEX13<='1' ; 
HEX14<='0' ; 
HEX15<='0' ; 
HEX16<='1' ;
		HEX20<='1' ; 
		HEX21<='0' ; 
		HEX22<='0' ; 
		HEX23<='0' ; 
		HEX24<='0' ; 
		HEX25<='0' ; 
		HEX26<='1' ;
HEX30<='0' ;
HEX31<='1' ;
HEX32<='0' ;
HEX33<='0' ;
HEX34<='0' ;
HEX35<='0' ;
HEX36<='1' ;
		HEX40<='1';
		HEX41<='1';
		HEX42<='1';
		HEX43<='1';
		HEX44<='1';
		HEX45<='1';
		HEX46<='1';
HEX50<='1';
HEX51<='1';
HEX52<='1';
HEX53<='1';
HEX54<='1';
HEX55<='1';
HEX56<='1';
		
	  i<="00100";
							--cas 5
	  when "00100" => 
	  HEX00<='1';
	  HEX01<='0';
	  HEX02<='0';	
	  HEX03<='1';
	  HEX04<='0';
	  HEX05<='0';
	  HEX06<='0' ;
HEX10<='1' ; 
HEX11<='1' ; 
HEX12<='1' ; 
HEX13<='0' ; 
HEX14<='0' ; 
HEX15<='0' ; 
HEX16<='1' ;	
		HEX20<='1' ; 
		HEX21<='1' ; 
		HEX22<='1' ; 
		HEX23<='1' ; 
		HEX24<='0' ; 
		HEX25<='0' ; 
		HEX26<='1' ;
HEX30<='1' ; 
HEX31<='0' ; 
HEX32<='0' ; 
HEX33<='0' ; 
HEX34<='0' ; 
HEX35<='0' ; 
HEX36<='1' ;
		HEX40<='0' ;
		HEX41<='1' ;
		HEX42<='0' ;
		HEX43<='0' ;
		HEX44<='0' ;
		HEX45<='0' ;
		HEX46<='1' ;
HEX50<='1';
HEX51<='1';
HEX52<='1';
HEX53<='1';
HEX54<='1';
HEX55<='1';
HEX56<='1';
		
	  i<="00101";
		when "00101" --cas 6
		=>
		HEX00<='0';
		HEX01<='1';
		HEX02<='1';
		HEX03<='0';
		HEX04<='0';
		HEX05<='0';
		HEX06<='0';
HEX10<='1' ; 
HEX11<='0' ; 
HEX12<='0' ; 
HEX13<='1' ; 
HEX14<='0' ; 
HEX15<='0' ; 
HEX16<='0' ;
			HEX20<='1' ; 
			HEX21<='1' ; 
			HEX22<='1' ; 
			HEX23<='0' ; 
			HEX24<='0' ; 
			HEX25<='0' ; 
			HEX26<='1' ;
HEX30<='1' ; 
HEX31<='1' ; 
HEX32<='1' ; 
HEX33<='1' ; 
HEX34<='0' ; 
HEX35<='0' ; 
HEX36<='1' ;
		HEX40<='1' ; 
		HEX41<='0' ; 
		HEX42<='0' ; 
		HEX43<='0' ; 
		HEX44<='0' ; 
		HEX45<='0' ; 
		HEX46<='1' ;
HEX50<='0' ;
HEX51<='1' ;
HEX52<='0' ;
HEX53<='0' ;
HEX54<='0' ;
HEX55<='0' ;
HEX56<='1' ;
	
		i<="00110";
		when "00110" --cas 7
		=>
		HEX00<='0';
		HEX01<='0';
		HEX02<='0';
		HEX03<='1';
		HEX04<='0';
		HEX05<='0';
		HEX06<='1';
HEX10<='0' ; 
HEX11<='1' ; 
HEX12<='1' ; 
HEX13<='0' ; 
HEX14<='0' ; 
HEX15<='0' ; 
HEX16<='0' ;
			HEX20<='1' ; 
			HEX21<='0' ; 
			HEX22<='0' ; 
			HEX23<='1' ; 
			HEX24<='0' ; 
			HEX25<='0' ; 
			HEX26<='0' ;
HEX30<='1' ; 
HEX31<='1' ; 
HEX32<='1' ; 
HEX33<='0' ; 
HEX34<='0' ; 
HEX35<='0' ; 
HEX36<='1' ;
		HEX40<='1' ; 
		HEX41<='1' ; 
		HEX42<='1' ; 
		HEX43<='1' ; 
		HEX44<='0' ; 
		HEX45<='0' ; 
		HEX46<='1' ;
HEX50<='1' ; 
HEX51<='0' ; 
HEX52<='0' ; 
HEX53<='0' ; 
HEX54<='0' ; 
HEX55<='0' ; 
HEX56<='1' ;
		
		i<="00111";
		when "00111" --cas 8
		=>
		HEX00<='1';
		HEX01<='1';
		HEX02<='1';
		HEX03<='1';
		HEX04<='1';
		HEX05<='1';
		HEX06<='1';
HEX10<='0' ; 
HEX11<='0' ; 
HEX12<='0' ; 
HEX13<='1' ; 
HEX14<='0' ; 
HEX15<='0' ; 
HEX16<='1' ;
			HEX20<='0' ; 
			HEX21<='1' ; 
			HEX22<='1' ; 
			HEX23<='0' ; 
			HEX24<='0' ; 
			HEX25<='0' ; 
			HEX26<='0' ;
HEX30<='1' ; 
HEX31<='0' ; 
HEX32<='0' ; 
HEX33<='1' ; 
HEX34<='0' ; 
HEX35<='0' ; 
HEX36<='0' ;
		HEX40<='1' ; 
		HEX41<='1' ; 
		HEX42<='1' ; 
		HEX43<='0' ; 
		HEX44<='0' ; 
		HEX45<='0' ; 
		HEX46<='1' ;
HEX50<='1' ; 
HEX51<='1' ; 
HEX52<='1' ; 
HEX53<='1' ; 
HEX54<='0' ; 
HEX55<='0' ; 
HEX56<='1' ;
		
		i<="01000";
		when "01000" --cas 9
		=>
		HEX00<='0';
		HEX01<='0';
		HEX02<='0';
		HEX03<='1';
		HEX04<='0';
		HEX05<='0';
		HEX06<='1';
HEX10<='1';
HEX11<='1';
HEX12<='1';
HEX13<='1';
HEX14<='1';
HEX15<='1';
HEX16<='1';
			HEX20<='0' ; 
			HEX21<='0' ; 
			HEX22<='0' ; 
			HEX23<='1' ; 
			HEX24<='0' ; 
			HEX25<='0' ; 
			HEX26<='1' ;
HEX30<='0' ; 
HEX31<='1' ; 
HEX32<='1' ; 
HEX33<='0' ; 
HEX34<='0' ; 
HEX35<='0' ; 
HEX36<='0' ;
		HEX40<='1' ; 
		HEX41<='0' ; 
		HEX42<='0' ; 
		HEX43<='1' ; 
		HEX44<='0' ; 
		HEX45<='0' ; 
		HEX46<='0' ;
HEX50<='1' ; 
HEX51<='1' ; 
HEX52<='1' ; 
HEX53<='0' ; 
HEX54<='0' ; 
HEX55<='0' ; 
HEX56<='1' ;
		
		i<="01001";
		when "01001" --cas 10
		=>
		HEX00<='0';
		HEX01<='0';
		HEX02<='0';
		HEX03<='1';
		HEX04<='0';
		HEX05<='0';
		HEX06<='0';
HEX10<='0' ; 
HEX11<='0' ; 
HEX12<='0' ; 
HEX13<='1' ; 
HEX14<='0' ; 
HEX15<='0' ; 
HEX16<='1' ;
			HEX20<='1';
			HEX21<='1';
			HEX22<='1';
			HEX23<='1';
			HEX24<='1';
			HEX25<='1';
			HEX26<='1';
HEX30<='0' ; 
HEX31<='0' ; 
HEX32<='0' ; 
HEX33<='1' ; 
HEX34<='0' ; 
HEX35<='0' ; 
HEX36<='1' ;
		HEX40<='0' ; 
		HEX41<='1' ; 
		HEX42<='1' ; 
		HEX43<='0' ; 
		HEX44<='0' ; 
		HEX45<='0' ; 
		HEX46<='0' ;
HEX50<='1' ; 
HEX51<='0' ; 
HEX52<='0' ; 
HEX53<='1' ; 
HEX54<='0' ; 
HEX55<='0' ; 
HEX56<='0' ;
		
		i<="01010";
		when "01010" --cas 11
		=>
		HEX00<='0';
		HEX01<='1';
		HEX02<='1';
		HEX03<='1';
		HEX04<='0';
		HEX05<='0';
		HEX06<='1';
HEX10<='0' ; 
HEX11<='0' ; 
HEX12<='0' ; 
HEX13<='1' ; 
HEX14<='0' ; 
HEX15<='0' ; 
HEX16<='0' ;
			HEX20<='0' ; 
			HEX21<='0' ; 
			HEX22<='0' ; 
			HEX23<='1' ; 
			HEX24<='0' ; 
			HEX25<='0' ; 
			HEX26<='1' ;
HEX30<='1';
HEX31<='1';
HEX32<='1';
HEX33<='1';
HEX34<='1';
HEX35<='1';
HEX36<='1';
		HEX40<='0' ; 
		HEX41<='0' ; 
		HEX42<='0' ; 
		HEX43<='1' ; 
		HEX44<='0' ; 
		HEX45<='0' ; 
		HEX46<='1' ;
HEX50<='0' ; 
HEX51<='1' ; 
HEX52<='1' ; 
HEX53<='0' ; 
HEX54<='0' ; 
HEX55<='0' ; 
HEX56<='0' ;
		
		i<="01011";
		when "01011" --cas 12
		=>
		HEX00<='0';
		HEX01<='1';
		HEX02<='1';
		HEX03<='1';
		HEX04<='0';
		HEX05<='0';
		HEX06<='1';
HEX10<='0' ; 
HEX11<='1' ; 
HEX12<='1' ; 
HEX13<='1' ; 
HEX14<='0' ; 
HEX15<='0' ; 
HEX16<='1' ;
			HEX20<='0' ; 
			HEX21<='0' ; 
			HEX22<='0' ; 
			HEX23<='1' ; 
			HEX24<='0' ; 
			HEX25<='0' ; 
			HEX26<='0' ;
HEX30<='0' ; 
HEX31<='0' ; 
HEX32<='0' ; 
HEX33<='1' ; 
HEX34<='0' ; 
HEX35<='0' ; 
HEX36<='1' ;
		HEX40<='1';
		HEX41<='1';
		HEX42<='1';
		HEX43<='1';
		HEX44<='1';
		HEX45<='1';
		HEX46<='1';
HEX50<='0' ; 
HEX51<='0' ; 
HEX52<='0' ; 
HEX53<='1' ; 
HEX54<='0' ; 
HEX55<='0' ; 
HEX56<='1' ;
		
		i<="01100";
		when "01100" --cas 13
		=>
		HEX00<='1';
		HEX01<='0';
		HEX02<='0';
		HEX03<='1';
		HEX04<='0';
		HEX05<='0';
		HEX06<='0';
HEX10<='0' ; 
HEX11<='1' ; 
HEX12<='1' ; 
HEX13<='1' ; 
HEX14<='0' ; 
HEX15<='0' ; 
HEX16<='1' ;
			HEX20<='0' ; 
			HEX21<='1' ; 
			HEX22<='1' ; 
			HEX23<='1' ; 
			HEX24<='0' ; 
			HEX25<='0' ; 
			HEX26<='1' ;
HEX30<='0' ; 
HEX31<='0' ; 
HEX32<='0' ; 
HEX33<='1' ; 
HEX34<='0' ; 
HEX35<='0' ; 
HEX36<='0' ;
		HEX40<='0' ; 
		HEX41<='0' ; 
		HEX42<='0' ; 
		HEX43<='1' ; 
		HEX44<='0' ; 
		HEX45<='0' ; 
		HEX46<='1' ;
HEX50<='1';
HEX51<='1';
HEX52<='1';
HEX53<='1';
HEX54<='1';
HEX55<='1';
HEX56<='1';
		
		i<="01101";
		when "01101" --cas 14
		=>
		HEX00<='1';
		HEX01<='1';
		HEX02<='1';
		HEX03<='1';
		HEX04<='0';
		HEX05<='0';
		HEX06<='1';
HEX10<='1' ; 
HEX11<='0' ; 
HEX12<='0' ; 
HEX13<='1' ; 
HEX14<='0' ; 
HEX15<='0' ; 
HEX16<='0' ;
			HEX20<='0' ; 
			HEX21<='1' ; 
			HEX22<='1' ; 
			HEX23<='1' ; 
			HEX24<='0' ; 
			HEX25<='0' ; 
			HEX26<='1' ;
HEX30<='0' ; 
HEX31<='1' ; 
HEX32<='1' ; 
HEX33<='1' ; 
HEX34<='0' ; 
HEX35<='0' ; 
HEX36<='1' ;
		HEX40<='0' ; 
		HEX41<='0' ; 
		HEX42<='0' ; 
		HEX43<='1' ; 
		HEX44<='0' ; 
		HEX45<='0' ; 
		HEX46<='0' ;
HEX50<='0' ; 
HEX51<='0' ; 
HEX52<='0' ; 
HEX53<='1' ; 
HEX54<='0' ; 
HEX55<='0' ; 
HEX56<='1' ;
	
		i<="01110";
		when "01110" --cas 15
		=>
		HEX00<='0';
		HEX01<='1';
		HEX02<='1';
		HEX03<='0';
		HEX04<='0';
		HEX05<='0';
		HEX06<='0';
HEX10<='1' ; 
HEX11<='1' ; 
HEX12<='1' ; 
HEX13<='1' ; 
HEX14<='0' ; 
HEX15<='0' ; 
HEX16<='1' ;
			HEX20<='1' ; 
			HEX21<='0' ; 
			HEX22<='0' ; 
			HEX23<='1' ; 
			HEX24<='0' ; 
			HEX25<='0' ; 
			HEX26<='0' ;
HEX30<='0' ; 
HEX31<='1' ; 
HEX32<='1' ; 
HEX33<='1' ; 
HEX34<='0' ; 
HEX35<='0' ; 
HEX36<='1' ;
		HEX40<='0' ; 
		HEX41<='1' ; 
		HEX42<='1' ; 
		HEX43<='1' ; 
		HEX44<='0' ; 
		HEX45<='0' ; 
		HEX46<='1' ;
HEX50<='0' ; 
HEX51<='0' ; 
HEX52<='0' ; 
HEX53<='1' ; 
HEX54<='0' ; 
HEX55<='0' ; 
HEX56<='0' ;
		
		i<="01111";
		when "01111" --cas 16
		=>
		HEX00<='1';
		HEX01<='0';
		HEX02<='0';
		HEX03<='0';
		HEX04<='0';
		HEX05<='0';
		HEX06<='1';
HEX10<='0' ; 
HEX11<='1' ; 
HEX12<='1' ; 
HEX13<='0' ; 
HEX14<='0' ; 
HEX15<='0' ; 
HEX16<='0' ;
			HEX20<='1' ; 
			HEX21<='1' ; 
			HEX22<='1' ; 
			HEX23<='1' ; 
			HEX24<='0' ; 
			HEX25<='0' ; 
			HEX26<='1' ;
HEX30<='1' ; 
HEX31<='0' ; 
HEX32<='0' ; 
HEX33<='1' ; 
HEX34<='0' ; 
HEX35<='0' ; 
HEX36<='0' ;
		HEX40<='0' ; 
		HEX41<='1' ; 
		HEX42<='1' ; 
		HEX43<='1' ; 
		HEX44<='0' ; 
		HEX45<='0' ; 
		HEX46<='1' ;
HEX50<='0' ; 
HEX51<='1' ; 
HEX52<='1' ; 
HEX53<='1' ; 
HEX54<='0' ; 
HEX55<='0' ; 
HEX56<='1' ;
		
		i<="10000";
		when "10000" --cas 17
		=>
		HEX00<='1';
		HEX01<='1';
		HEX02<='1';
		HEX03<='1';
		HEX04<='1';
		HEX05<='1';
		HEX06<='1';
HEX10<='1' ; 
HEX11<='0' ; 
HEX12<='0' ; 
HEX13<='0' ; 
HEX14<='0' ; 
HEX15<='0' ; 
HEX16<='1' ;
			HEX20<='0' ; 
			HEX21<='1' ; 
			HEX22<='1' ; 
			HEX23<='0' ; 
			HEX24<='0' ; 
			HEX25<='0' ; 
			HEX26<='0' ;
HEX30<='1' ; 
HEX31<='1' ; 
HEX32<='1' ; 
HEX33<='1' ; 
HEX34<='0' ; 
HEX35<='0' ; 
HEX36<='1' ;
		HEX40<='1' ; 
		HEX41<='0' ; 
		HEX42<='0' ; 
		HEX43<='1' ; 
		HEX44<='0' ; 
		HEX45<='0' ; 
		HEX46<='0' ;
HEX50<='0' ; 
HEX51<='1' ; 
HEX52<='1' ; 
HEX53<='1' ; 
HEX54<='0' ; 
HEX55<='0' ; 
HEX56<='1' ;
		
		i<="10001";
		when "10001" --cas 18
		=>
		HEX00<='1';
		HEX01<='1';
		HEX02<='1';
		HEX03<='1';
		HEX04<='1';
		HEX05<='1';
		HEX06<='1';
HEX10<='1';
HEX11<='1';
HEX12<='1';
HEX13<='1';
HEX14<='1';
HEX15<='1';
HEX16<='1';
			HEX20<='1' ; 
			HEX21<='0' ; 
			HEX22<='0' ; 
			HEX23<='0' ; 
			HEX24<='0' ; 
			HEX25<='0' ; 
			HEX26<='1' ;
HEX30<='0' ; 
HEX31<='1' ; 
HEX32<='1' ; 
HEX33<='0' ; 
HEX34<='0' ; 
HEX35<='0' ; 
HEX36<='0' ;
		HEX40<='1' ; 
		HEX41<='1' ; 
		HEX42<='1' ; 
		HEX43<='1' ; 
		HEX44<='0' ; 
		HEX45<='0' ; 
		HEX46<='1' ;
HEX50<='1' ; 
HEX51<='0' ; 
HEX52<='0' ; 
HEX53<='1' ; 
HEX54<='0' ; 
HEX55<='0' ; 
HEX56<='0' ;
		
		i<="10010";
		when "10010" --cas 19
		=>
		HEX00<='1';
		HEX01<='1';
		HEX02<='1';
		HEX03<='1';
		HEX04<='1';
		HEX05<='1';
		HEX06<='1';
HEX10<='1';
HEX11<='1';
HEX12<='1';
HEX13<='1';
HEX14<='1';
HEX15<='1';
HEX16<='1';
			HEX20<='1';
			HEX21<='1';
			HEX22<='1';
			HEX23<='1';
			HEX24<='1';
			HEX25<='1';
			HEX26<='1';
HEX30<='1' ; 
HEX31<='0' ; 
HEX32<='0' ; 
HEX33<='0' ; 
HEX34<='0' ; 
HEX35<='0' ; 
HEX36<='1' ;
		HEX40<='0' ; 
		HEX41<='1' ; 
		HEX42<='1' ; 
		HEX43<='0' ; 
		HEX44<='0' ; 
		HEX45<='0' ; 
		HEX46<='0' ;
HEX50<='1' ; 
HEX51<='1' ; 
HEX52<='1' ; 
HEX53<='1' ; 
HEX54<='0' ; 
HEX55<='0' ; 
HEX56<='1' ;
		
		i<="10011";
		when "10011" --cas 20
		=>
		HEX00<='1';
		HEX01<='1';
		HEX02<='1';
		HEX03<='1';
		HEX04<='1';
		HEX05<='1';
		HEX06<='1';
HEX10<='1';
HEX11<='1';
HEX12<='1';
HEX13<='1';
HEX14<='1';
HEX15<='1';
HEX16<='1';
			HEX20<='1';
			HEX21<='1';
			HEX22<='1';
			HEX23<='1';
			HEX24<='1';
			HEX25<='1';
			HEX26<='1';
HEX30<='1';
HEX31<='1';
HEX32<='1';
HEX33<='1';
HEX34<='1';
HEX35<='1';
HEX36<='1';
		HEX40<='1' ; 
		HEX41<='0' ; 
		HEX42<='0' ; 
		HEX43<='0' ; 
		HEX44<='0' ; 
		HEX45<='0' ; 
		HEX46<='1' ;
HEX50<='0' ; 
HEX51<='1' ; 
HEX52<='1' ; 
HEX53<='0' ; 
HEX54<='0' ; 
HEX55<='0' ; 
HEX56<='0' ;
		
		i<="10100";
		when "10100" --cas 21
		=>
		HEX00<='1';
		HEX01<='1';
		HEX02<='1';
		HEX03<='1';
		HEX04<='1';
		HEX05<='1';
		HEX06<='1';
HEX10<='1';
HEX11<='1';
HEX12<='1';
HEX13<='1';
HEX14<='1';
HEX15<='1';
HEX16<='1';
			HEX20<='1';
			HEX21<='1';
			HEX22<='1';
			HEX23<='1';
			HEX24<='1';
			HEX25<='1';
			HEX26<='1';
HEX30<='1';
HEX31<='1';
HEX32<='1';
HEX33<='1';
HEX34<='1';
HEX35<='1';
HEX36<='1';
		HEX40<='1' ; 
		HEX41<='1' ; 
		HEX42<='1' ; 
		HEX43<='1' ; 
		HEX44<='1' ; 
		HEX45<='1' ; 
		HEX46<='1' ;
HEX50<='1' ; 
HEX51<='0' ; 
HEX52<='0' ; 
HEX53<='0' ; 
HEX54<='0' ; 
HEX55<='0' ; 
HEX56<='1' ;
		
		i<="10101";
		when "10101" --cas 22
		=>
		HEX00<='1';
		HEX01<='1';
		HEX02<='1';
		HEX03<='1';
		HEX04<='1';
		HEX05<='1';
		HEX06<='1';
HEX10<='1';
HEX11<='1';
HEX12<='1';
HEX13<='1';
HEX14<='1';
HEX15<='1';
HEX16<='1';
			HEX20<='1';
			HEX21<='1';
			HEX22<='1';
			HEX23<='1';
			HEX24<='1';
			HEX25<='1';
			HEX26<='1';
HEX30<='1';
HEX31<='1';
HEX32<='1';
HEX33<='1';
HEX34<='1';
HEX35<='1';
HEX36<='1';
		HEX40<='1' ; 
		HEX41<='1' ; 
		HEX42<='1' ; 
		HEX43<='1' ; 
		HEX44<='1' ; 
		HEX45<='1' ; 
		HEX46<='1' ;
HEX50<='1' ; 
HEX51<='1' ; 
HEX52<='1' ; 
HEX53<='1' ; 
HEX54<='1' ; 
HEX55<='1' ; 
HEX56<='1' ;
		
		i<="10110";
		when "10110" --cas 23
		=>
		HEX00<='1';
		HEX01<='1';
		HEX02<='1';
		HEX03<='1';
		HEX04<='1';
		HEX05<='1';
		HEX06<='1';
HEX10<='1';
HEX11<='1';
HEX12<='1';
HEX13<='1';
HEX14<='1';
HEX15<='1';
HEX16<='1';
			HEX20<='1';
			HEX21<='1';
			HEX22<='1';
			HEX23<='1';
			HEX24<='1';
			HEX25<='1';
			HEX26<='1';
HEX30<='1';
HEX31<='1';
HEX32<='1';
HEX33<='1';
HEX34<='1';
HEX35<='1';
HEX36<='1';
		HEX40<='1' ; 
		HEX41<='1' ; 
		HEX42<='1' ; 
		HEX43<='1' ; 
		HEX44<='1' ; 
		HEX45<='1' ; 
		HEX46<='1' ;
HEX50<='1' ; 
HEX51<='1' ; 
HEX52<='1' ; 
HEX53<='1' ; 
HEX54<='1' ; 
HEX55<='1' ; 
HEX56<='1' ;
		
		i<="00000";

		
		when others =>
	  
	  i<="00000";
		end case;
		
	end if; 
	if(SW0='0') then 
	case i is  
		when "00000" => 
								--cas 1	
	  HEX00 <= '0';
	  HEX01 <= '1';
	  HEX02 <= '0';
	  HEX03 <= '0';
	  HEX04 <= '0';
	  HEX05 <= '0';
	  HEX06 <= '1';
HEX10<='1';
HEX11<='1';
HEX12<='1';
HEX13<='1';
HEX14<='1';
HEX15<='1';
HEX16<='1';
			HEX20<='1';
			HEX21<='1';
			HEX22<='1';
			HEX23<='1';
			HEX24<='1';
			HEX25<='1';
			HEX26<='1';
HEX30<='1';
HEX31<='1';
HEX32<='1';
HEX33<='1';
HEX34<='1';
HEX35<='1';
HEX36<='1';	
		HEX40<='1';
		HEX41<='1';
		HEX42<='1';
		HEX43<='1';
		HEX44<='1';
		HEX45<='1';
		HEX46<='1';
HEX50<='1';
HEX51<='1';
HEX52<='1';
HEX53<='1';
HEX54<='1';
HEX55<='1';
HEX56<='1';
	
	  
	  
								--cas 2
	  when "00001" => 
	  HEX00<='1';
	  HEX01<='0';
	  HEX02<='0';
	  HEX03<='0';
	  HEX04<='0';
	  HEX05<='0';
	  HEX06<='1' ;
HEX10<='0' ;
HEX11<='1' ;
HEX12<='0' ;
HEX13<='0' ;
HEX14<='0' ;
HEX15<='0' ;
HEX16<='1' ;
		HEX20<='1';
		HEX21<='1';
		HEX22<='1';
		HEX23<='1';
		HEX24<='1';
		HEX25<='1';
		HEX26<='1';
HEX30<='1';
HEX31<='1';
HEX32<='1';
HEX33<='1';
HEX34<='1';
HEX35<='1';
HEX36<='1';
		HEX40<='1';
		HEX41<='1';
		HEX42<='1';
		HEX43<='1';
		HEX44<='1';
		HEX45<='1';
		HEX46<='1';
HEX50<='1';
HEX51<='1';
HEX52<='1';
HEX53<='1';
HEX54<='1';
HEX55<='1';
HEX56<='1';
		

								--cas 3
	  when "00010" => 
	  HEX00<='1';
	  HEX01<='1';
	  HEX02<='1';
	  HEX03<='1';
	  HEX04<='0';
	  HEX05<='0';
	  HEX06<='1' ;
HEX10<='1' ; 
HEX11<='0' ; 
HEX12<='0' ; 
HEX13<='0' ; 
HEX14<='0' ; 
HEX15<='0' ; 
HEX16<='1' ;
		HEX20<='0' ;
		HEX21<='1' ;
		HEX22<='0' ;
		HEX23<='0' ;
		HEX24<='0' ;
		HEX25<='0' ;
		HEX26<='1' ;
HEX30<='1';
HEX31<='1';
HEX32<='1';
HEX33<='1';
HEX34<='1';
HEX35<='1';
HEX36<='1';
		HEX40<='1';
		HEX41<='1';
		HEX42<='1';
		HEX43<='1';
		HEX44<='1';
		HEX45<='1';
		HEX46<='1';
HEX50<='1';
HEX51<='1';
HEX52<='1';
HEX53<='1';
HEX54<='1';
HEX55<='1';
HEX56<='1';
		
							--cas 4
	  when "00011" => 
	  HEX00<='1';
	  HEX01<='1';
	  HEX02<='1';
	  HEX03<='0';
	  HEX04<='0';
	  HEX05<='0';
	  HEX06<='1' ;
HEX10<='1' ; 
HEX11<='1' ; 
HEX12<='1' ; 
HEX13<='1' ; 
HEX14<='0' ; 
HEX15<='0' ; 
HEX16<='1' ;
		HEX20<='1' ; 
		HEX21<='0' ; 
		HEX22<='0' ; 
		HEX23<='0' ; 
		HEX24<='0' ; 
		HEX25<='0' ; 
		HEX26<='1' ;
HEX30<='0' ;
HEX31<='1' ;
HEX32<='0' ;
HEX33<='0' ;
HEX34<='0' ;
HEX35<='0' ;
HEX36<='1' ;
		HEX40<='1';
		HEX41<='1';
		HEX42<='1';
		HEX43<='1';
		HEX44<='1';
		HEX45<='1';
		HEX46<='1';
HEX50<='1';
HEX51<='1';
HEX52<='1';
HEX53<='1';
HEX54<='1';
HEX55<='1';
HEX56<='1';
		
							--cas 5
	  when "00100" => 
	  HEX00<='1';
	  HEX01<='0';
	  HEX02<='0';	
	  HEX03<='1';
	  HEX04<='0';
	  HEX05<='0';
	  HEX06<='0' ;
HEX10<='1' ; 
HEX11<='1' ; 
HEX12<='1' ; 
HEX13<='0' ; 
HEX14<='0' ; 
HEX15<='0' ; 
HEX16<='1' ;	
		HEX20<='1' ; 
		HEX21<='1' ; 
		HEX22<='1' ; 
		HEX23<='1' ; 
		HEX24<='0' ; 
		HEX25<='0' ; 
		HEX26<='1' ;
HEX30<='1' ; 
HEX31<='0' ; 
HEX32<='0' ; 
HEX33<='0' ; 
HEX34<='0' ; 
HEX35<='0' ; 
HEX36<='1' ;
		HEX40<='0' ;
		HEX41<='1' ;
		HEX42<='0' ;
		HEX43<='0' ;
		HEX44<='0' ;
		HEX45<='0' ;
		HEX46<='1' ;
HEX50<='1';
HEX51<='1';
HEX52<='1';
HEX53<='1';
HEX54<='1';
HEX55<='1';
HEX56<='1';
		
		when "00101" --cas 6
		=>
		HEX00<='0';
		HEX01<='1';
		HEX02<='1';
		HEX03<='0';
		HEX04<='0';
		HEX05<='0';
		HEX06<='0';
HEX10<='1' ; 
HEX11<='0' ; 
HEX12<='0' ; 
HEX13<='1' ; 
HEX14<='0' ; 
HEX15<='0' ; 
HEX16<='0' ;
			HEX20<='1' ; 
			HEX21<='1' ; 
			HEX22<='1' ; 
			HEX23<='0' ; 
			HEX24<='0' ; 
			HEX25<='0' ; 
			HEX26<='1' ;
HEX30<='1' ; 
HEX31<='1' ; 
HEX32<='1' ; 
HEX33<='1' ; 
HEX34<='0' ; 
HEX35<='0' ; 
HEX36<='1' ;
		HEX40<='1' ; 
		HEX41<='0' ; 
		HEX42<='0' ; 
		HEX43<='0' ; 
		HEX44<='0' ; 
		HEX45<='0' ; 
		HEX46<='1' ;
HEX50<='0' ;
HEX51<='1' ;
HEX52<='0' ;
HEX53<='0' ;
HEX54<='0' ;
HEX55<='0' ;
HEX56<='1' ;
	
		when "00110" --cas 7
		=>
		HEX00<='0';
		HEX01<='0';
		HEX02<='0';
		HEX03<='1';
		HEX04<='0';
		HEX05<='0';
		HEX06<='1';
HEX10<='0' ; 
HEX11<='1' ; 
HEX12<='1' ; 
HEX13<='0' ; 
HEX14<='0' ; 
HEX15<='0' ; 
HEX16<='0' ;
			HEX20<='1' ; 
			HEX21<='0' ; 
			HEX22<='0' ; 
			HEX23<='1' ; 
			HEX24<='0' ; 
			HEX25<='0' ; 
			HEX26<='0' ;
HEX30<='1' ; 
HEX31<='1' ; 
HEX32<='1' ; 
HEX33<='0' ; 
HEX34<='0' ; 
HEX35<='0' ; 
HEX36<='1' ;
		HEX40<='1' ; 
		HEX41<='1' ; 
		HEX42<='1' ; 
		HEX43<='1' ; 
		HEX44<='0' ; 
		HEX45<='0' ; 
		HEX46<='1' ;
HEX50<='1' ; 
HEX51<='0' ; 
HEX52<='0' ; 
HEX53<='0' ; 
HEX54<='0' ; 
HEX55<='0' ; 
HEX56<='1' ;
		
		when "00111" --cas 8
		=>
		HEX00<='1';
		HEX01<='1';
		HEX02<='1';
		HEX03<='1';
		HEX04<='1';
		HEX05<='1';
		HEX06<='1';
HEX10<='0' ; 
HEX11<='0' ; 
HEX12<='0' ; 
HEX13<='1' ; 
HEX14<='0' ; 
HEX15<='0' ; 
HEX16<='1' ;
			HEX20<='0' ; 
			HEX21<='1' ; 
			HEX22<='1' ; 
			HEX23<='0' ; 
			HEX24<='0' ; 
			HEX25<='0' ; 
			HEX26<='0' ;
HEX30<='1' ; 
HEX31<='0' ; 
HEX32<='0' ; 
HEX33<='1' ; 
HEX34<='0' ; 
HEX35<='0' ; 
HEX36<='0' ;
		HEX40<='1' ; 
		HEX41<='1' ; 
		HEX42<='1' ; 
		HEX43<='0' ; 
		HEX44<='0' ; 
		HEX45<='0' ; 
		HEX46<='1' ;
HEX50<='1' ; 
HEX51<='1' ; 
HEX52<='1' ; 
HEX53<='1' ; 
HEX54<='0' ; 
HEX55<='0' ; 
HEX56<='1' ;
		
		when "01000" --cas 9
		=>
		HEX00<='0';
		HEX01<='0';
		HEX02<='0';
		HEX03<='1';
		HEX04<='0';
		HEX05<='0';
		HEX06<='1';
HEX10<='1';
HEX11<='1';
HEX12<='1';
HEX13<='1';
HEX14<='1';
HEX15<='1';
HEX16<='1';
			HEX20<='0' ; 
			HEX21<='0' ; 
			HEX22<='0' ; 
			HEX23<='1' ; 
			HEX24<='0' ; 
			HEX25<='0' ; 
			HEX26<='1' ;
HEX30<='0' ; 
HEX31<='1' ; 
HEX32<='1' ; 
HEX33<='0' ; 
HEX34<='0' ; 
HEX35<='0' ; 
HEX36<='0' ;
		HEX40<='1' ; 
		HEX41<='0' ; 
		HEX42<='0' ; 
		HEX43<='1' ; 
		HEX44<='0' ; 
		HEX45<='0' ; 
		HEX46<='0' ;
HEX50<='1' ; 
HEX51<='1' ; 
HEX52<='1' ; 
HEX53<='0' ; 
HEX54<='0' ; 
HEX55<='0' ; 
HEX56<='1' ;
		
		when "01001" --cas 10
		=>
		HEX00<='0';
		HEX01<='0';
		HEX02<='0';
		HEX03<='1';
		HEX04<='0';
		HEX05<='0';
		HEX06<='0';
HEX10<='0' ; 
HEX11<='0' ; 
HEX12<='0' ; 
HEX13<='1' ; 
HEX14<='0' ; 
HEX15<='0' ; 
HEX16<='1' ;
			HEX20<='1';
			HEX21<='1';
			HEX22<='1';
			HEX23<='1';
			HEX24<='1';
			HEX25<='1';
			HEX26<='1';
HEX30<='0' ; 
HEX31<='0' ; 
HEX32<='0' ; 
HEX33<='1' ; 
HEX34<='0' ; 
HEX35<='0' ; 
HEX36<='1' ;
		HEX40<='0' ; 
		HEX41<='1' ; 
		HEX42<='1' ; 
		HEX43<='0' ; 
		HEX44<='0' ; 
		HEX45<='0' ; 
		HEX46<='0' ;
HEX50<='1' ; 
HEX51<='0' ; 
HEX52<='0' ; 
HEX53<='1' ; 
HEX54<='0' ; 
HEX55<='0' ; 
HEX56<='0' ;
		when "01010" --cas 11
		=>
		HEX00<='0';
		HEX01<='1';
		HEX02<='1';
		HEX03<='1';
		HEX04<='0';
		HEX05<='0';
		HEX06<='1';
HEX10<='0' ; 
HEX11<='0' ; 
HEX12<='0' ; 
HEX13<='1' ; 
HEX14<='0' ; 
HEX15<='0' ; 
HEX16<='0' ;
			HEX20<='0' ; 
			HEX21<='0' ; 
			HEX22<='0' ; 
			HEX23<='1' ; 
			HEX24<='0' ; 
			HEX25<='0' ; 
			HEX26<='1' ;
HEX30<='1';
HEX31<='1';
HEX32<='1';
HEX33<='1';
HEX34<='1';
HEX35<='1';
HEX36<='1';
		HEX40<='0' ; 
		HEX41<='0' ; 
		HEX42<='0' ; 
		HEX43<='1' ; 
		HEX44<='0' ; 
		HEX45<='0' ; 
		HEX46<='1' ;
HEX50<='0' ; 
HEX51<='1' ; 
HEX52<='1' ; 
HEX53<='0' ; 
HEX54<='0' ; 
HEX55<='0' ; 
HEX56<='0' ;
		
		when "01011" --cas 12
		=>
		HEX00<='0';
		HEX01<='1';
		HEX02<='1';
		HEX03<='1';
		HEX04<='0';
		HEX05<='0';
		HEX06<='1';
HEX10<='0' ; 
HEX11<='1' ; 
HEX12<='1' ; 
HEX13<='1' ; 
HEX14<='0' ; 
HEX15<='0' ; 
HEX16<='1' ;
			HEX20<='0' ; 
			HEX21<='0' ; 
			HEX22<='0' ; 
			HEX23<='1' ; 
			HEX24<='0' ; 
			HEX25<='0' ; 
			HEX26<='0' ;
HEX30<='0' ; 
HEX31<='0' ; 
HEX32<='0' ; 
HEX33<='1' ; 
HEX34<='0' ; 
HEX35<='0' ; 
HEX36<='1' ;
		HEX40<='1';
		HEX41<='1';
		HEX42<='1';
		HEX43<='1';
		HEX44<='1';
		HEX45<='1';
		HEX46<='1';
HEX50<='0' ; 
HEX51<='0' ; 
HEX52<='0' ; 
HEX53<='1' ; 
HEX54<='0' ; 
HEX55<='0' ; 
HEX56<='1' ;
		
		when "01100" --cas 13
		=>
		HEX00<='1';
		HEX01<='0';
		HEX02<='0';
		HEX03<='1';
		HEX04<='0';
		HEX05<='0';
		HEX06<='0';
HEX10<='0' ; 
HEX11<='1' ; 
HEX12<='1' ; 
HEX13<='1' ; 
HEX14<='0' ; 
HEX15<='0' ; 
HEX16<='1' ;
			HEX20<='0' ; 
			HEX21<='1' ; 
			HEX22<='1' ; 
			HEX23<='1' ; 
			HEX24<='0' ; 
			HEX25<='0' ; 
			HEX26<='1' ;
HEX30<='0' ; 
HEX31<='0' ; 
HEX32<='0' ; 
HEX33<='1' ; 
HEX34<='0' ; 
HEX35<='0' ; 
HEX36<='0' ;
		HEX40<='0' ; 
		HEX41<='0' ; 
		HEX42<='0' ; 
		HEX43<='1' ; 
		HEX44<='0' ; 
		HEX45<='0' ; 
		HEX46<='1' ;
HEX50<='1';
HEX51<='1';
HEX52<='1';
HEX53<='1';
HEX54<='1';
HEX55<='1';
HEX56<='1';
		
		
		when "01101" --cas 14
		=>
		HEX00<='1';
		HEX01<='1';
		HEX02<='1';
		HEX03<='1';
		HEX04<='0';
		HEX05<='0';
		HEX06<='1';
HEX10<='1' ; 
HEX11<='0' ; 
HEX12<='0' ; 
HEX13<='1' ; 
HEX14<='0' ; 
HEX15<='0' ; 
HEX16<='0' ;
			HEX20<='0' ; 
			HEX21<='1' ; 
			HEX22<='1' ; 
			HEX23<='1' ; 
			HEX24<='0' ; 
			HEX25<='0' ; 
			HEX26<='1' ;
HEX30<='0' ; 
HEX31<='1' ; 
HEX32<='1' ; 
HEX33<='1' ; 
HEX34<='0' ; 
HEX35<='0' ; 
HEX36<='1' ;
		HEX40<='0' ; 
		HEX41<='0' ; 
		HEX42<='0' ; 
		HEX43<='1' ; 
		HEX44<='0' ; 
		HEX45<='0' ; 
		HEX46<='0' ;
HEX50<='0' ; 
HEX51<='0' ; 
HEX52<='0' ; 
HEX53<='1' ; 
HEX54<='0' ; 
HEX55<='0' ; 
HEX56<='1' ;
	
		when "01110" --cas 15
		=>
		HEX00<='0';
		HEX01<='1';
		HEX02<='1';
		HEX03<='0';
		HEX04<='0';
		HEX05<='0';
		HEX06<='0';
HEX10<='1' ; 
HEX11<='1' ; 
HEX12<='1' ; 
HEX13<='1' ; 
HEX14<='0' ; 
HEX15<='0' ; 
HEX16<='1' ;
			HEX20<='1' ; 
			HEX21<='0' ; 
			HEX22<='0' ; 
			HEX23<='1' ; 
			HEX24<='0' ; 
			HEX25<='0' ; 
			HEX26<='0' ;
HEX30<='0' ; 
HEX31<='1' ; 
HEX32<='1' ; 
HEX33<='1' ; 
HEX34<='0' ; 
HEX35<='0' ; 
HEX36<='1' ;
		HEX40<='0' ; 
		HEX41<='1' ; 
		HEX42<='1' ; 
		HEX43<='1' ; 
		HEX44<='0' ; 
		HEX45<='0' ; 
		HEX46<='1' ;
HEX50<='0' ; 
HEX51<='0' ; 
HEX52<='0' ; 
HEX53<='1' ; 
HEX54<='0' ; 
HEX55<='0' ; 
HEX56<='0' ;
		
		
		when "01111" --cas 16
		=>
		HEX00<='1';
		HEX01<='0';
		HEX02<='0';
		HEX03<='0';
		HEX04<='0';
		HEX05<='0';
		HEX06<='1';
HEX10<='0' ; 
HEX11<='1' ; 
HEX12<='1' ; 
HEX13<='0' ; 
HEX14<='0' ; 
HEX15<='0' ; 
HEX16<='0' ;
			HEX20<='1' ; 
			HEX21<='1' ; 
			HEX22<='1' ; 
			HEX23<='1' ; 
			HEX24<='0' ; 
			HEX25<='0' ; 
			HEX26<='1' ;
HEX30<='1' ; 
HEX31<='0' ; 
HEX32<='0' ; 
HEX33<='1' ; 
HEX34<='0' ; 
HEX35<='0' ; 
HEX36<='0' ;
		HEX40<='0' ; 
		HEX41<='1' ; 
		HEX42<='1' ; 
		HEX43<='1' ; 
		HEX44<='0' ; 
		HEX45<='0' ; 
		HEX46<='1' ;
HEX50<='0' ; 
HEX51<='1' ; 
HEX52<='1' ; 
HEX53<='1' ; 
HEX54<='0' ; 
HEX55<='0' ; 
HEX56<='1' ;
		
		
		when "10000" --cas 17
		=>
		HEX00<='1';
		HEX01<='1';
		HEX02<='1';
		HEX03<='1';
		HEX04<='1';
		HEX05<='1';
		HEX06<='1';
HEX10<='1' ; 
HEX11<='0' ; 
HEX12<='0' ; 
HEX13<='0' ; 
HEX14<='0' ; 
HEX15<='0' ; 
HEX16<='1' ;
			HEX20<='0' ; 
			HEX21<='1' ; 
			HEX22<='1' ; 
			HEX23<='0' ; 
			HEX24<='0' ; 
			HEX25<='0' ; 
			HEX26<='0' ;
HEX30<='1' ; 
HEX31<='1' ; 
HEX32<='1' ; 
HEX33<='1' ; 
HEX34<='0' ; 
HEX35<='0' ; 
HEX36<='1' ;
		HEX40<='1' ; 
		HEX41<='0' ; 
		HEX42<='0' ; 
		HEX43<='1' ; 
		HEX44<='0' ; 
		HEX45<='0' ; 
		HEX46<='0' ;
HEX50<='0' ; 
HEX51<='1' ; 
HEX52<='1' ; 
HEX53<='1' ; 
HEX54<='0' ; 
HEX55<='0' ; 
HEX56<='1' ;
		
		
		when "10001" --cas 18
		=>
		HEX00<='1';
		HEX01<='1';
		HEX02<='1';
		HEX03<='1';
		HEX04<='1';
		HEX05<='1';
		HEX06<='1';
HEX10<='1';
HEX11<='1';
HEX12<='1';
HEX13<='1';
HEX14<='1';
HEX15<='1';
HEX16<='1';
			HEX20<='1' ; 
			HEX21<='0' ; 
			HEX22<='0' ; 
			HEX23<='0' ; 
			HEX24<='0' ; 
			HEX25<='0' ; 
			HEX26<='1' ;
HEX30<='0' ; 
HEX31<='1' ; 
HEX32<='1' ; 
HEX33<='0' ; 
HEX34<='0' ; 
HEX35<='0' ; 
HEX36<='0' ;
		HEX40<='1' ; 
		HEX41<='1' ; 
		HEX42<='1' ; 
		HEX43<='1' ; 
		HEX44<='0' ; 
		HEX45<='0' ; 
		HEX46<='1' ;
HEX50<='1' ; 
HEX51<='0' ; 
HEX52<='0' ; 
HEX53<='1' ; 
HEX54<='0' ; 
HEX55<='0' ; 
HEX56<='0' ;
	
		when "10010" --cas 19
		=>
		HEX00<='1';
		HEX01<='1';
		HEX02<='1';
		HEX03<='1';
		HEX04<='1';
		HEX05<='1';
		HEX06<='1';
HEX10<='1';
HEX11<='1';
HEX12<='1';
HEX13<='1';
HEX14<='1';
HEX15<='1';
HEX16<='1';
			HEX20<='1';
			HEX21<='1';
			HEX22<='1';
			HEX23<='1';
			HEX24<='1';
			HEX25<='1';
			HEX26<='1';
HEX30<='1' ; 
HEX31<='0' ; 
HEX32<='0' ; 
HEX33<='0' ; 
HEX34<='0' ; 
HEX35<='0' ; 
HEX36<='1' ;
		HEX40<='0' ; 
		HEX41<='1' ; 
		HEX42<='1' ; 
		HEX43<='0' ; 
		HEX44<='0' ; 
		HEX45<='0' ; 
		HEX46<='0' ;
HEX50<='1' ; 
HEX51<='1' ; 
HEX52<='1' ; 
HEX53<='1' ; 
HEX54<='0' ; 
HEX55<='0' ; 
HEX56<='1' ;
		
		
		when "10011" --cas 20
		=>
		HEX00<='1';
		HEX01<='1';
		HEX02<='1';
		HEX03<='1';
		HEX04<='1';
		HEX05<='1';
		HEX06<='1';
HEX10<='1';
HEX11<='1';
HEX12<='1';
HEX13<='1';
HEX14<='1';
HEX15<='1';
HEX16<='1';
			HEX20<='1';
			HEX21<='1';
			HEX22<='1';
			HEX23<='1';
			HEX24<='1';
			HEX25<='1';
			HEX26<='1';
HEX30<='1';
HEX31<='1';
HEX32<='1';
HEX33<='1';
HEX34<='1';
HEX35<='1';
HEX36<='1';
		HEX40<='1' ; 
		HEX41<='0' ; 
		HEX42<='0' ; 
		HEX43<='0' ; 
		HEX44<='0' ; 
		HEX45<='0' ; 
		HEX46<='1' ;
HEX50<='0' ; 
HEX51<='1' ; 
HEX52<='1' ; 
HEX53<='0' ; 
HEX54<='0' ; 
HEX55<='0' ; 
HEX56<='0' ;
		
		
		when "10100" --cas 21
		=>
		HEX00<='1';
		HEX01<='1';
		HEX02<='1';
		HEX03<='1';
		HEX04<='1';
		HEX05<='1';
		HEX06<='1';
HEX10<='1';
HEX11<='1';
HEX12<='1';
HEX13<='1';
HEX14<='1';
HEX15<='1';
HEX16<='1';
			HEX20<='1';
			HEX21<='1';
			HEX22<='1';
			HEX23<='1';
			HEX24<='1';
			HEX25<='1';
			HEX26<='1';
HEX30<='1';
HEX31<='1';
HEX32<='1';
HEX33<='1';
HEX34<='1';
HEX35<='1';
HEX36<='1';
		HEX40<='1' ; 
		HEX41<='1' ; 
		HEX42<='1' ; 
		HEX43<='1' ; 
		HEX44<='1' ; 
		HEX45<='1' ; 
		HEX46<='1' ;
HEX50<='1' ; 
HEX51<='0' ; 
HEX52<='0' ; 
HEX53<='0' ; 
HEX54<='0' ; 
HEX55<='0' ; 
HEX56<='1' ;
		
		
		when "10101" --cas 22
		=>
		HEX00<='1';
		HEX01<='1';
		HEX02<='1';
		HEX03<='1';
		HEX04<='1';
		HEX05<='1';
		HEX06<='1';
HEX10<='1';
HEX11<='1';
HEX12<='1';
HEX13<='1';
HEX14<='1';
HEX15<='1';
HEX16<='1';
			HEX20<='1';
			HEX21<='1';
			HEX22<='1';
			HEX23<='1';
			HEX24<='1';
			HEX25<='1';
			HEX26<='1';
HEX30<='1';
HEX31<='1';
HEX32<='1';
HEX33<='1';
HEX34<='1';
HEX35<='1';
HEX36<='1';
		HEX40<='1' ; 
		HEX41<='1' ; 
		HEX42<='1' ; 
		HEX43<='1' ; 
		HEX44<='1' ; 
		HEX45<='1' ; 
		HEX46<='1' ;
HEX50<='1' ; 
HEX51<='1' ; 
HEX52<='1' ; 
HEX53<='1' ; 
HEX54<='1' ; 
HEX55<='1' ; 
HEX56<='1' ;
		
		
		when "10110" --cas 23
		=>
		HEX00<='1';
		HEX01<='1';
		HEX02<='1';
		HEX03<='1';
		HEX04<='1';
		HEX05<='1';
		HEX06<='1';
HEX10<='1';
HEX11<='1';
HEX12<='1';
HEX13<='1';
HEX14<='1';
HEX15<='1';
HEX16<='1';
			HEX20<='1';
			HEX21<='1';
			HEX22<='1';
			HEX23<='1';
			HEX24<='1';
			HEX25<='1';
			HEX26<='1';
HEX30<='1';
HEX31<='1';
HEX32<='1';
HEX33<='1';
HEX34<='1';
HEX35<='1';
HEX36<='1';
		HEX40<='1' ; 
		HEX41<='1' ; 
		HEX42<='1' ; 
		HEX43<='1' ; 
		HEX44<='1' ; 
		HEX45<='1' ; 
		HEX46<='1' ;
HEX50<='1' ; 
HEX51<='1' ; 
HEX52<='1' ; 
HEX53<='1' ; 
HEX54<='1' ; 
HEX55<='1' ; 
HEX56<='1' ;
		
		

		
		when others =>
	  
	  i<="00000";
		end case;
	
		end if;
		if(sw1='0') then 
		case i is  
		when "00000" => 
								--cas 1	
	  HEX00 <= '0';
	  HEX01 <= '1';
	  HEX02 <= '0';
	  HEX03 <= '0';
	  HEX04 <= '0';
	  HEX05 <= '0';
	  HEX06 <= '1';
HEX10<='1';
HEX11<='1';
HEX12<='1';
HEX13<='1';
HEX14<='1';
HEX15<='1';
HEX16<='1';
			HEX20<='1';
			HEX21<='1';
			HEX22<='1';
			HEX23<='1';
			HEX24<='1';
			HEX25<='1';
			HEX26<='1';
HEX30<='1';
HEX31<='1';
HEX32<='1';
HEX33<='1';
HEX34<='1';
HEX35<='1';
HEX36<='1';	
		HEX40<='1';
		HEX41<='1';
		HEX42<='1';
		HEX43<='1';
		HEX44<='1';
		HEX45<='1';
		HEX46<='1';
HEX50<='1';
HEX51<='1';
HEX52<='1';
HEX53<='1';
HEX54<='1';
HEX55<='1';
HEX56<='1';
	
	  
	  i <= "10110";
	  
								--cas 2
	  when "00001" => 
	  HEX00<='1';
	  HEX01<='0';
	  HEX02<='0';
	  HEX03<='0';
	  HEX04<='0';
	  HEX05<='0';
	  HEX06<='1' ;
HEX10<='0' ;
HEX11<='1' ;
HEX12<='0' ;
HEX13<='0' ;
HEX14<='0' ;
HEX15<='0' ;
HEX16<='1' ;
		HEX20<='1';
		HEX21<='1';
		HEX22<='1';
		HEX23<='1';
		HEX24<='1';
		HEX25<='1';
		HEX26<='1';
HEX30<='1';
HEX31<='1';
HEX32<='1';
HEX33<='1';
HEX34<='1';
HEX35<='1';
HEX36<='1';
		HEX40<='1';
		HEX41<='1';
		HEX42<='1';
		HEX43<='1';
		HEX44<='1';
		HEX45<='1';
		HEX46<='1';
HEX50<='1';
HEX51<='1';
HEX52<='1';
HEX53<='1';
HEX54<='1';
HEX55<='1';
HEX56<='1';
		

	  i<="00000";
								--cas 3
	  when "00010" => 
	  HEX00<='1';
	  HEX01<='1';
	  HEX02<='1';
	  HEX03<='1';
	  HEX04<='0';
	  HEX05<='0';
	  HEX06<='1' ;
HEX10<='1' ; 
HEX11<='0' ; 
HEX12<='0' ; 
HEX13<='0' ; 
HEX14<='0' ; 
HEX15<='0' ; 
HEX16<='1' ;
		HEX20<='0' ;
		HEX21<='1' ;
		HEX22<='0' ;
		HEX23<='0' ;
		HEX24<='0' ;
		HEX25<='0' ;
		HEX26<='1' ;
HEX30<='1';
HEX31<='1';
HEX32<='1';
HEX33<='1';
HEX34<='1';
HEX35<='1';
HEX36<='1';
		HEX40<='1';
		HEX41<='1';
		HEX42<='1';
		HEX43<='1';
		HEX44<='1';
		HEX45<='1';
		HEX46<='1';
HEX50<='1';
HEX51<='1';
HEX52<='1';
HEX53<='1';
HEX54<='1';
HEX55<='1';
HEX56<='1';
		
	  i<="00001";
							--cas 4
	  when "00011" => 
	  HEX00<='1';
	  HEX01<='1';
	  HEX02<='1';
	  HEX03<='0';
	  HEX04<='0';
	  HEX05<='0';
	  HEX06<='1' ;
HEX10<='1' ; 
HEX11<='1' ; 
HEX12<='1' ; 
HEX13<='1' ; 
HEX14<='0' ; 
HEX15<='0' ; 
HEX16<='1' ;
		HEX20<='1' ; 
		HEX21<='0' ; 
		HEX22<='0' ; 
		HEX23<='0' ; 
		HEX24<='0' ; 
		HEX25<='0' ; 
		HEX26<='1' ;
HEX30<='0' ;
HEX31<='1' ;
HEX32<='0' ;
HEX33<='0' ;
HEX34<='0' ;
HEX35<='0' ;
HEX36<='1' ;
		HEX40<='1';
		HEX41<='1';
		HEX42<='1';
		HEX43<='1';
		HEX44<='1';
		HEX45<='1';
		HEX46<='1';
HEX50<='1';
HEX51<='1';
HEX52<='1';
HEX53<='1';
HEX54<='1';
HEX55<='1';
HEX56<='1';
		
	  i<="00010";
							--cas 5
	  when "00100" => 
	  HEX00<='1';
	  HEX01<='0';
	  HEX02<='0';	
	  HEX03<='1';
	  HEX04<='0';
	  HEX05<='0';
	  HEX06<='0' ;
HEX10<='1' ; 
HEX11<='1' ; 
HEX12<='1' ; 
HEX13<='0' ; 
HEX14<='0' ; 
HEX15<='0' ; 
HEX16<='1' ;	
		HEX20<='1' ; 
		HEX21<='1' ; 
		HEX22<='1' ; 
		HEX23<='1' ; 
		HEX24<='0' ; 
		HEX25<='0' ; 
		HEX26<='1' ;
HEX30<='1' ; 
HEX31<='0' ; 
HEX32<='0' ; 
HEX33<='0' ; 
HEX34<='0' ; 
HEX35<='0' ; 
HEX36<='1' ;
		HEX40<='0' ;
		HEX41<='1' ;
		HEX42<='0' ;
		HEX43<='0' ;
		HEX44<='0' ;
		HEX45<='0' ;
		HEX46<='1' ;
HEX50<='1';
HEX51<='1';
HEX52<='1';
HEX53<='1';
HEX54<='1';
HEX55<='1';
HEX56<='1';
		
	  i<="00011";
		when "00101" --cas 6
		=>
		HEX00<='0';
		HEX01<='1';
		HEX02<='1';
		HEX03<='0';
		HEX04<='0';
		HEX05<='0';
		HEX06<='0';
HEX10<='1' ; 
HEX11<='0' ; 
HEX12<='0' ; 
HEX13<='1' ; 
HEX14<='0' ; 
HEX15<='0' ; 
HEX16<='0' ;
			HEX20<='1' ; 
			HEX21<='1' ; 
			HEX22<='1' ; 
			HEX23<='0' ; 
			HEX24<='0' ; 
			HEX25<='0' ; 
			HEX26<='1' ;
HEX30<='1' ; 
HEX31<='1' ; 
HEX32<='1' ; 
HEX33<='1' ; 
HEX34<='0' ; 
HEX35<='0' ; 
HEX36<='1' ;
		HEX40<='1' ; 
		HEX41<='0' ; 
		HEX42<='0' ; 
		HEX43<='0' ; 
		HEX44<='0' ; 
		HEX45<='0' ; 
		HEX46<='1' ;
HEX50<='0' ;
HEX51<='1' ;
HEX52<='0' ;
HEX53<='0' ;
HEX54<='0' ;
HEX55<='0' ;
HEX56<='1' ;
	
		i<="00100";
		when "00110" --cas 7
		=>
		HEX00<='0';
		HEX01<='0';
		HEX02<='0';
		HEX03<='1';
		HEX04<='0';
		HEX05<='0';
		HEX06<='1';
HEX10<='0' ; 
HEX11<='1' ; 
HEX12<='1' ; 
HEX13<='0' ; 
HEX14<='0' ; 
HEX15<='0' ; 
HEX16<='0' ;
			HEX20<='1' ; 
			HEX21<='0' ; 
			HEX22<='0' ; 
			HEX23<='1' ; 
			HEX24<='0' ; 
			HEX25<='0' ; 
			HEX26<='0' ;
HEX30<='1' ; 
HEX31<='1' ; 
HEX32<='1' ; 
HEX33<='0' ; 
HEX34<='0' ; 
HEX35<='0' ; 
HEX36<='1' ;
		HEX40<='1' ; 
		HEX41<='1' ; 
		HEX42<='1' ; 
		HEX43<='1' ; 
		HEX44<='0' ; 
		HEX45<='0' ; 
		HEX46<='1' ;
HEX50<='1' ; 
HEX51<='0' ; 
HEX52<='0' ; 
HEX53<='0' ; 
HEX54<='0' ; 
HEX55<='0' ; 
HEX56<='1' ;
		
		i<="00101";
		when "00111" --cas 8
		=>
		HEX00<='1';
		HEX01<='1';
		HEX02<='1';
		HEX03<='1';
		HEX04<='1';
		HEX05<='1';
		HEX06<='1';
HEX10<='0' ; 
HEX11<='0' ; 
HEX12<='0' ; 
HEX13<='1' ; 
HEX14<='0' ; 
HEX15<='0' ; 
HEX16<='1' ;
			HEX20<='0' ; 
			HEX21<='1' ; 
			HEX22<='1' ; 
			HEX23<='0' ; 
			HEX24<='0' ; 
			HEX25<='0' ; 
			HEX26<='0' ;
HEX30<='1' ; 
HEX31<='0' ; 
HEX32<='0' ; 
HEX33<='1' ; 
HEX34<='0' ; 
HEX35<='0' ; 
HEX36<='0' ;
		HEX40<='1' ; 
		HEX41<='1' ; 
		HEX42<='1' ; 
		HEX43<='0' ; 
		HEX44<='0' ; 
		HEX45<='0' ; 
		HEX46<='1' ;
HEX50<='1' ; 
HEX51<='1' ; 
HEX52<='1' ; 
HEX53<='1' ; 
HEX54<='0' ; 
HEX55<='0' ; 
HEX56<='1' ;
		
		i<="00110";
		when "01000" --cas 9
		=>
		HEX00<='0';
		HEX01<='0';
		HEX02<='0';
		HEX03<='1';
		HEX04<='0';
		HEX05<='0';
		HEX06<='1';
HEX10<='1';
HEX11<='1';
HEX12<='1';
HEX13<='1';
HEX14<='1';
HEX15<='1';
HEX16<='1';
			HEX20<='0' ; 
			HEX21<='0' ; 
			HEX22<='0' ; 
			HEX23<='1' ; 
			HEX24<='0' ; 
			HEX25<='0' ; 
			HEX26<='1' ;
HEX30<='0' ; 
HEX31<='1' ; 
HEX32<='1' ; 
HEX33<='0' ; 
HEX34<='0' ; 
HEX35<='0' ; 
HEX36<='0' ;
		HEX40<='1' ; 
		HEX41<='0' ; 
		HEX42<='0' ; 
		HEX43<='1' ; 
		HEX44<='0' ; 
		HEX45<='0' ; 
		HEX46<='0' ;
HEX50<='1' ; 
HEX51<='1' ; 
HEX52<='1' ; 
HEX53<='0' ; 
HEX54<='0' ; 
HEX55<='0' ; 
HEX56<='1' ;
		
		i<="00111";
		when "01001" --cas 10
		=>
		HEX00<='0';
		HEX01<='0';
		HEX02<='0';
		HEX03<='1';
		HEX04<='0';
		HEX05<='0';
		HEX06<='0';
HEX10<='0' ; 
HEX11<='0' ; 
HEX12<='0' ; 
HEX13<='1' ; 
HEX14<='0' ; 
HEX15<='0' ; 
HEX16<='1' ;
			HEX20<='1';
			HEX21<='1';
			HEX22<='1';
			HEX23<='1';
			HEX24<='1';
			HEX25<='1';
			HEX26<='1';
HEX30<='0' ; 
HEX31<='0' ; 
HEX32<='0' ; 
HEX33<='1' ; 
HEX34<='0' ; 
HEX35<='0' ; 
HEX36<='1' ;
		HEX40<='0' ; 
		HEX41<='1' ; 
		HEX42<='1' ; 
		HEX43<='0' ; 
		HEX44<='0' ; 
		HEX45<='0' ; 
		HEX46<='0' ;
HEX50<='1' ; 
HEX51<='0' ; 
HEX52<='0' ; 
HEX53<='1' ; 
HEX54<='0' ; 
HEX55<='0' ; 
HEX56<='0' ;
		
		i<="01000";
		when "01010" --cas 11
		=>
		HEX00<='0';
		HEX01<='1';
		HEX02<='1';
		HEX03<='1';
		HEX04<='0';
		HEX05<='0';
		HEX06<='1';
HEX10<='0' ; 
HEX11<='0' ; 
HEX12<='0' ; 
HEX13<='1' ; 
HEX14<='0' ; 
HEX15<='0' ; 
HEX16<='0' ;
			HEX20<='0' ; 
			HEX21<='0' ; 
			HEX22<='0' ; 
			HEX23<='1' ; 
			HEX24<='0' ; 
			HEX25<='0' ; 
			HEX26<='1' ;
HEX30<='1';
HEX31<='1';
HEX32<='1';
HEX33<='1';
HEX34<='1';
HEX35<='1';
HEX36<='1';
		HEX40<='0' ; 
		HEX41<='0' ; 
		HEX42<='0' ; 
		HEX43<='1' ; 
		HEX44<='0' ; 
		HEX45<='0' ; 
		HEX46<='1' ;
HEX50<='0' ; 
HEX51<='1' ; 
HEX52<='1' ; 
HEX53<='0' ; 
HEX54<='0' ; 
HEX55<='0' ; 
HEX56<='0' ;
		
		i<="01001";
		when "01011" --cas 12
		=>
		HEX00<='0';
		HEX01<='1';
		HEX02<='1';
		HEX03<='1';
		HEX04<='0';
		HEX05<='0';
		HEX06<='1';
HEX10<='0' ; 
HEX11<='1' ; 
HEX12<='1' ; 
HEX13<='1' ; 
HEX14<='0' ; 
HEX15<='0' ; 
HEX16<='1' ;
			HEX20<='0' ; 
			HEX21<='0' ; 
			HEX22<='0' ; 
			HEX23<='1' ; 
			HEX24<='0' ; 
			HEX25<='0' ; 
			HEX26<='0' ;
HEX30<='0' ; 
HEX31<='0' ; 
HEX32<='0' ; 
HEX33<='1' ; 
HEX34<='0' ; 
HEX35<='0' ; 
HEX36<='1' ;
		HEX40<='1';
		HEX41<='1';
		HEX42<='1';
		HEX43<='1';
		HEX44<='1';
		HEX45<='1';
		HEX46<='1';
HEX50<='0' ; 
HEX51<='0' ; 
HEX52<='0' ; 
HEX53<='1' ; 
HEX54<='0' ; 
HEX55<='0' ; 
HEX56<='1' ;
		
		i<="01010";
		when "01100" --cas 13
		=>
		HEX00<='1';
		HEX01<='0';
		HEX02<='0';
		HEX03<='1';
		HEX04<='0';
		HEX05<='0';
		HEX06<='0';
HEX10<='0' ; 
HEX11<='1' ; 
HEX12<='1' ; 
HEX13<='1' ; 
HEX14<='0' ; 
HEX15<='0' ; 
HEX16<='1' ;
			HEX20<='0' ; 
			HEX21<='1' ; 
			HEX22<='1' ; 
			HEX23<='1' ; 
			HEX24<='0' ; 
			HEX25<='0' ; 
			HEX26<='1' ;
HEX30<='0' ; 
HEX31<='0' ; 
HEX32<='0' ; 
HEX33<='1' ; 
HEX34<='0' ; 
HEX35<='0' ; 
HEX36<='0' ;
		HEX40<='0' ; 
		HEX41<='0' ; 
		HEX42<='0' ; 
		HEX43<='1' ; 
		HEX44<='0' ; 
		HEX45<='0' ; 
		HEX46<='1' ;
HEX50<='1';
HEX51<='1';
HEX52<='1';
HEX53<='1';
HEX54<='1';
HEX55<='1';
HEX56<='1';
		
		i<="01011";
		when "01101" --cas 14
		=>
		HEX00<='1';
		HEX01<='1';
		HEX02<='1';
		HEX03<='1';
		HEX04<='0';
		HEX05<='0';
		HEX06<='1';
HEX10<='1' ; 
HEX11<='0' ; 
HEX12<='0' ; 
HEX13<='1' ; 
HEX14<='0' ; 
HEX15<='0' ; 
HEX16<='0' ;
			HEX20<='0' ; 
			HEX21<='1' ; 
			HEX22<='1' ; 
			HEX23<='1' ; 
			HEX24<='0' ; 
			HEX25<='0' ; 
			HEX26<='1' ;
HEX30<='0' ; 
HEX31<='1' ; 
HEX32<='1' ; 
HEX33<='1' ; 
HEX34<='0' ; 
HEX35<='0' ; 
HEX36<='1' ;
		HEX40<='0' ; 
		HEX41<='0' ; 
		HEX42<='0' ; 
		HEX43<='1' ; 
		HEX44<='0' ; 
		HEX45<='0' ; 
		HEX46<='0' ;
HEX50<='0' ; 
HEX51<='0' ; 
HEX52<='0' ; 
HEX53<='1' ; 
HEX54<='0' ; 
HEX55<='0' ; 
HEX56<='1' ;
	
		i<="01100";
		when "01110" --cas 15
		=>
		HEX00<='0';
		HEX01<='1';
		HEX02<='1';
		HEX03<='0';
		HEX04<='0';
		HEX05<='0';
		HEX06<='0';
HEX10<='1' ; 
HEX11<='1' ; 
HEX12<='1' ; 
HEX13<='1' ; 
HEX14<='0' ; 
HEX15<='0' ; 
HEX16<='1' ;
			HEX20<='1' ; 
			HEX21<='0' ; 
			HEX22<='0' ; 
			HEX23<='1' ; 
			HEX24<='0' ; 
			HEX25<='0' ; 
			HEX26<='0' ;
HEX30<='0' ; 
HEX31<='1' ; 
HEX32<='1' ; 
HEX33<='1' ; 
HEX34<='0' ; 
HEX35<='0' ; 
HEX36<='1' ;
		HEX40<='0' ; 
		HEX41<='1' ; 
		HEX42<='1' ; 
		HEX43<='1' ; 
		HEX44<='0' ; 
		HEX45<='0' ; 
		HEX46<='1' ;
HEX50<='0' ; 
HEX51<='0' ; 
HEX52<='0' ; 
HEX53<='1' ; 
HEX54<='0' ; 
HEX55<='0' ; 
HEX56<='0' ;
		
		i<="01101";
		when "01111" --cas 16
		=>
		HEX00<='1';
		HEX01<='0';
		HEX02<='0';
		HEX03<='0';
		HEX04<='0';
		HEX05<='0';
		HEX06<='1';
HEX10<='0' ; 
HEX11<='1' ; 
HEX12<='1' ; 
HEX13<='0' ; 
HEX14<='0' ; 
HEX15<='0' ; 
HEX16<='0' ;
			HEX20<='1' ; 
			HEX21<='1' ; 
			HEX22<='1' ; 
			HEX23<='1' ; 
			HEX24<='0' ; 
			HEX25<='0' ; 
			HEX26<='1' ;
HEX30<='1' ; 
HEX31<='0' ; 
HEX32<='0' ; 
HEX33<='1' ; 
HEX34<='0' ; 
HEX35<='0' ; 
HEX36<='0' ;
		HEX40<='0' ; 
		HEX41<='1' ; 
		HEX42<='1' ; 
		HEX43<='1' ; 
		HEX44<='0' ; 
		HEX45<='0' ; 
		HEX46<='1' ;
HEX50<='0' ; 
HEX51<='1' ; 
HEX52<='1' ; 
HEX53<='1' ; 
HEX54<='0' ; 
HEX55<='0' ; 
HEX56<='1' ;
		
		i<="01110";
		when "10000" --cas 17
		=>
		HEX00<='1';
		HEX01<='1';
		HEX02<='1';
		HEX03<='1';
		HEX04<='1';
		HEX05<='1';
		HEX06<='1';
HEX10<='1' ; 
HEX11<='0' ; 
HEX12<='0' ; 
HEX13<='0' ; 
HEX14<='0' ; 
HEX15<='0' ; 
HEX16<='1' ;
			HEX20<='0' ; 
			HEX21<='1' ; 
			HEX22<='1' ; 
			HEX23<='0' ; 
			HEX24<='0' ; 
			HEX25<='0' ; 
			HEX26<='0' ;
HEX30<='1' ; 
HEX31<='1' ; 
HEX32<='1' ; 
HEX33<='1' ; 
HEX34<='0' ; 
HEX35<='0' ; 
HEX36<='1' ;
		HEX40<='1' ; 
		HEX41<='0' ; 
		HEX42<='0' ; 
		HEX43<='1' ; 
		HEX44<='0' ; 
		HEX45<='0' ; 
		HEX46<='0' ;
HEX50<='0' ; 
HEX51<='1' ; 
HEX52<='1' ; 
HEX53<='1' ; 
HEX54<='0' ; 
HEX55<='0' ; 
HEX56<='1' ;
		
		i<="01111";
		when "10001" --cas 18
		=>
		HEX00<='1';
		HEX01<='1';
		HEX02<='1';
		HEX03<='1';
		HEX04<='1';
		HEX05<='1';
		HEX06<='1';
HEX10<='1';
HEX11<='1';
HEX12<='1';
HEX13<='1';
HEX14<='1';
HEX15<='1';
HEX16<='1';
			HEX20<='1' ; 
			HEX21<='0' ; 
			HEX22<='0' ; 
			HEX23<='0' ; 
			HEX24<='0' ; 
			HEX25<='0' ; 
			HEX26<='1' ;
HEX30<='0' ; 
HEX31<='1' ; 
HEX32<='1' ; 
HEX33<='0' ; 
HEX34<='0' ; 
HEX35<='0' ; 
HEX36<='0' ;
		HEX40<='1' ; 
		HEX41<='1' ; 
		HEX42<='1' ; 
		HEX43<='1' ; 
		HEX44<='0' ; 
		HEX45<='0' ; 
		HEX46<='1' ;
HEX50<='1' ; 
HEX51<='0' ; 
HEX52<='0' ; 
HEX53<='1' ; 
HEX54<='0' ; 
HEX55<='0' ; 
HEX56<='0' ;
		
		i<="10000";
		when "10010" --cas 19
		=>
		HEX00<='1';
		HEX01<='1';
		HEX02<='1';
		HEX03<='1';
		HEX04<='1';
		HEX05<='1';
		HEX06<='1';
HEX10<='1';
HEX11<='1';
HEX12<='1';
HEX13<='1';
HEX14<='1';
HEX15<='1';
HEX16<='1';
			HEX20<='1';
			HEX21<='1';
			HEX22<='1';
			HEX23<='1';
			HEX24<='1';
			HEX25<='1';
			HEX26<='1';
HEX30<='1' ; 
HEX31<='0' ; 
HEX32<='0' ; 
HEX33<='0' ; 
HEX34<='0' ; 
HEX35<='0' ; 
HEX36<='1' ;
		HEX40<='0' ; 
		HEX41<='1' ; 
		HEX42<='1' ; 
		HEX43<='0' ; 
		HEX44<='0' ; 
		HEX45<='0' ; 
		HEX46<='0' ;
HEX50<='1' ; 
HEX51<='1' ; 
HEX52<='1' ; 
HEX53<='1' ; 
HEX54<='0' ; 
HEX55<='0' ; 
HEX56<='1' ;
		
		i<="10001";
		when "10011" --cas 20
		=>
		HEX00<='1';
		HEX01<='1';
		HEX02<='1';
		HEX03<='1';
		HEX04<='1';
		HEX05<='1';
		HEX06<='1';
HEX10<='1';
HEX11<='1';
HEX12<='1';
HEX13<='1';
HEX14<='1';
HEX15<='1';
HEX16<='1';
			HEX20<='1';
			HEX21<='1';
			HEX22<='1';
			HEX23<='1';
			HEX24<='1';
			HEX25<='1';
			HEX26<='1';
HEX30<='1';
HEX31<='1';
HEX32<='1';
HEX33<='1';
HEX34<='1';
HEX35<='1';
HEX36<='1';
		HEX40<='1' ; 
		HEX41<='0' ; 
		HEX42<='0' ; 
		HEX43<='0' ; 
		HEX44<='0' ; 
		HEX45<='0' ; 
		HEX46<='1' ;
HEX50<='0' ; 
HEX51<='1' ; 
HEX52<='1' ; 
HEX53<='0' ; 
HEX54<='0' ; 
HEX55<='0' ; 
HEX56<='0' ;
		
		i<="10010";
		when "10100" --cas 21
		=>
		HEX00<='1';
		HEX01<='1';
		HEX02<='1';
		HEX03<='1';
		HEX04<='1';
		HEX05<='1';
		HEX06<='1';
HEX10<='1';
HEX11<='1';
HEX12<='1';
HEX13<='1';
HEX14<='1';
HEX15<='1';
HEX16<='1';
			HEX20<='1';
			HEX21<='1';
			HEX22<='1';
			HEX23<='1';
			HEX24<='1';
			HEX25<='1';
			HEX26<='1';
HEX30<='1';
HEX31<='1';
HEX32<='1';
HEX33<='1';
HEX34<='1';
HEX35<='1';
HEX36<='1';
		HEX40<='1' ; 
		HEX41<='1' ; 
		HEX42<='1' ; 
		HEX43<='1' ; 
		HEX44<='1' ; 
		HEX45<='1' ; 
		HEX46<='1' ;
HEX50<='1' ; 
HEX51<='0' ; 
HEX52<='0' ; 
HEX53<='0' ; 
HEX54<='0' ; 
HEX55<='0' ; 
HEX56<='1' ;
		
		i<="10011";
		when "10101" --cas 22
		=>
		HEX00<='1';
		HEX01<='1';
		HEX02<='1';
		HEX03<='1';
		HEX04<='1';
		HEX05<='1';
		HEX06<='1';
HEX10<='1';
HEX11<='1';
HEX12<='1';
HEX13<='1';
HEX14<='1';
HEX15<='1';
HEX16<='1';
			HEX20<='1';
			HEX21<='1';
			HEX22<='1';
			HEX23<='1';
			HEX24<='1';
			HEX25<='1';
			HEX26<='1';
HEX30<='1';
HEX31<='1';
HEX32<='1';
HEX33<='1';
HEX34<='1';
HEX35<='1';
HEX36<='1';
		HEX40<='1' ; 
		HEX41<='1' ; 
		HEX42<='1' ; 
		HEX43<='1' ; 
		HEX44<='1' ; 
		HEX45<='1' ; 
		HEX46<='1' ;
HEX50<='1' ; 
HEX51<='1' ; 
HEX52<='1' ; 
HEX53<='1' ; 
HEX54<='1' ; 
HEX55<='1' ; 
HEX56<='1' ;
		
		i<="10100";
		when "10110" --cas 23
		=>
		HEX00<='1';
		HEX01<='1';
		HEX02<='1';
		HEX03<='1';
		HEX04<='1';
		HEX05<='1';
		HEX06<='1';
HEX10<='1';
HEX11<='1';
HEX12<='1';
HEX13<='1';
HEX14<='1';
HEX15<='1';
HEX16<='1';
			HEX20<='1';
			HEX21<='1';
			HEX22<='1';
			HEX23<='1';
			HEX24<='1';
			HEX25<='1';
			HEX26<='1';
HEX30<='1';
HEX31<='1';
HEX32<='1';
HEX33<='1';
HEX34<='1';
HEX35<='1';
HEX36<='1';
		HEX40<='1' ; 
		HEX41<='1' ; 
		HEX42<='1' ; 
		HEX43<='1' ; 
		HEX44<='1' ; 
		HEX45<='1' ; 
		HEX46<='1' ;
HEX50<='1' ; 
HEX51<='1' ; 
HEX52<='1' ; 
HEX53<='1' ; 
HEX54<='1' ; 
HEX55<='1' ; 
HEX56<='1' ;
		
		i<="10101";

		
		when others =>
	  
	  i<="00000";
		end case;
		end if;
 end if;
end process;
END behavioral;
